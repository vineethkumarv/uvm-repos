module one;
initial begin
  $display("hi");
end 
endmodule
